`timescale 1 ns / 1 ps

module ander (a, b, result);

    input a,b;
    output result;

    assign result = a & b;

endmodule
