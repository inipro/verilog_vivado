��f u n c t i o n   [ 1 5 : 0 ]   m u l t i p l y _ f u n c ;  
         i n p u t   [ 7 : 0 ]   a , b ;  
         r e g   [ 1 5 : 0 ]   c ;    
 b e g i n  
         c   =   a   *   b ;  
         m u l t i p l y _ f u n c   =   c ;  
 e n d  
 e n d f u n c t i o n  
 �  
 t a s k   m u l t i p l y _ t a s k ;  
         i n p u t   [ 7 : 0 ]   a , b ;  
         o u t p u t   [ 1 5 : 0 ]   c ;    
 b e g i n  
         c   =   a   *   b ;    
 e n d  
 e n d t a s k  
 